package fir_coeffs_pkg;
    localparam int N = 102;

    // Floating-point coefficients (double precision)
    const real COEFFS_FLOAT [0:N-1] = '{
        -0.0002346183,
        -0.0008799227,
        -0.0023164192,
        -0.0049397725,
        -0.0090752608,
        -0.0148083095,
        -0.0218158808,
        -0.0292573076,
        -0.0357908499,
        -0.0397601007,
        -0.0395483907,
        -0.0340378651,
        -0.0230543059,
        -0.0076493289,
        0.0099110385,
        0.0265162461,
        0.0388980676,
        0.0444812470,
        0.0421601395,
        0.0327487395,
        0.0189157430,
        0.0045595494,
        -0.0062461700,
        -0.0104473244,
        -0.0069751998,
        0.0028484929,
        0.0156480166,
        0.0270182290,
        0.0329482535,
        0.0311939240,
        0.0221277947,
        0.0087376308,
        -0.0042874202,
        -0.0121316481,
        -0.0115850856,
        -0.0023336911,
        0.0126856588,
        0.0280717799,
        0.0377110577,
        0.0369657987,
        0.0245747778,
        0.0035798330,
        -0.0191304328,
        -0.0346333259,
        -0.0346565754,
        -0.0143270413,
        0.0258994195,
        0.0797986251,
        0.1366591724,
        0.1839794519,
        0.2108194094,
        0.2108194094,
        0.1839794519,
        0.1366591724,
        0.0797986251,
        0.0258994195,
        -0.0143270413,
        -0.0346565754,
        -0.0346333259,
        -0.0191304328,
        0.0035798330,
        0.0245747778,
        0.0369657987,
        0.0377110577,
        0.0280717799,
        0.0126856588,
        -0.0023336911,
        -0.0115850856,
        -0.0121316481,
        -0.0042874202,
        0.0087376308,
        0.0221277947,
        0.0311939240,
        0.0329482535,
        0.0270182290,
        0.0156480166,
        0.0028484929,
        -0.0069751998,
        -0.0104473244,
        -0.0062461700,
        0.0045595494,
        0.0189157430,
        0.0327487395,
        0.0421601395,
        0.0444812470,
        0.0388980676,
        0.0265162461,
        0.0099110385,
        -0.0076493289,
        -0.0230543059,
        -0.0340378651,
        -0.0395483907,
        -0.0397601007,
        -0.0357908499,
        -0.0292573076,
        -0.0218158808,
        -0.0148083095,
        -0.0090752608,
        -0.0049397725,
        -0.0023164192,
        -0.0008799227,
        -0.0002346183
    };

    // Fixed-point coefficients (Q15 format)
    const logic signed [15:0] COEFFS_FIXED [0:N-1] = '{
        -16'sd8,
        -16'sd29,
        -16'sd76,
        -16'sd162,
        -16'sd297,
        -16'sd485,
        -16'sd715,
        -16'sd959,
        -16'sd1173,
        -16'sd1303,
        -16'sd1296,
        -16'sd1115,
        -16'sd755,
        -16'sd251,
        16'sd325,
        16'sd869,
        16'sd1275,
        16'sd1458,
        16'sd1382,
        16'sd1073,
        16'sd620,
        16'sd149,
        -16'sd205,
        -16'sd342,
        -16'sd229,
        16'sd93,
        16'sd513,
        16'sd885,
        16'sd1080,
        16'sd1022,
        16'sd725,
        16'sd286,
        -16'sd140,
        -16'sd398,
        -16'sd380,
        -16'sd76,
        16'sd416,
        16'sd920,
        16'sd1236,
        16'sd1211,
        16'sd805,
        16'sd117,
        -16'sd627,
        -16'sd1135,
        -16'sd1136,
        -16'sd469,
        16'sd849,
        16'sd2615,
        16'sd4478,
        16'sd6029,
        16'sd6908,
        16'sd6908,
        16'sd6029,
        16'sd4478,
        16'sd2615,
        16'sd849,
        -16'sd469,
        -16'sd1136,
        -16'sd1135,
        -16'sd627,
        16'sd117,
        16'sd805,
        16'sd1211,
        16'sd1236,
        16'sd920,
        16'sd416,
        -16'sd76,
        -16'sd380,
        -16'sd398,
        -16'sd140,
        16'sd286,
        16'sd725,
        16'sd1022,
        16'sd1080,
        16'sd885,
        16'sd513,
        16'sd93,
        -16'sd229,
        -16'sd342,
        -16'sd205,
        16'sd149,
        16'sd620,
        16'sd1073,
        16'sd1382,
        16'sd1458,
        16'sd1275,
        16'sd869,
        16'sd325,
        -16'sd251,
        -16'sd755,
        -16'sd1115,
        -16'sd1296,
        -16'sd1303,
        -16'sd1173,
        -16'sd959,
        -16'sd715,
        -16'sd485,
        -16'sd297,
        -16'sd162,
        -16'sd76,
        -16'sd29,
        -16'sd8
    };
endpackage
